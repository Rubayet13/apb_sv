package env_pkg;
        import agent_pkg::*;
        `include "apb_scb.sv"
        `include "apb_env.sv"
endpackage 