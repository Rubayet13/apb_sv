package agent_pkg;

    `include "apb_trans.sv"
    `include "apb_driver.sv"
    `include "apb_generator.sv"
    `include "apb_monitor.sv"

endpackage 
